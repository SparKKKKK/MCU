module fetch();
input 
output

